*
* OPAMP MACRO MODEL (INTERMEDIATE LEVEL)
*
*                IN+ IN- OUT  VCC  VEE
*.SUBCKT OPAMP    1   2   81   101   102 
* Change order to match spice opamp pins 1-5   
*                IN+ IN- VCC   VEE  OUT
.SUBCKT OPAMP    1   2   101   102  81 
Q1	5 1	7	NPN
Q2	6 2	8	NPN
RC1	101	5	95.49
RC2	101	6	95.49
RE1	7	4	43.79
RE2	8	4	43.79
I1	4	102	0.001
*
* OPEN-LOOP GAIN, FIRST POLE AND SLEW RATE
G1	100 10	6 5 0.0104719
RP1	10	100	9.549MEG
CP1	10	100	0.0016667UF
*
*OUTPUT STAGE
EOUT	80 100	10 100	1
RO	80	81	100
*
* INTERNAL REFERENCE
RREF1	101	103	100K
RREF2	103	102	100K
EREF	100 0	103 0 1
R100	100	0	1MEG
*
.model NPN  NPN(BF=50000)
*

.print v(1)

.ENDS
