* Schematic : /home/lroot/Desktop/sedra-spice/ex5.1.4/nmos-id-vds-char.sch
* Component Definitions
M1 1 2 0 0 nmos_enhancement_mosfet l=10u w=400u
Vds 1 0 DC 10V
Vgs 2 0 DC 5V

* Model Definitions
.MODEL nmos_enhancement_mosfet NMOS (kp=20u Vto=+2 lambda=0)

* NG-Spice Simulation Commands
*.DC Vds 0v 10v 100mv
*.PRINT DC I(Vds) V(1)

.control

echo ++++++++++++++++++++++++++++++++++
echo Starting of control section

let loopLet = 0
set loopSet = 0
foreach lmb 0 0.05 0.1
  * we could have just done "let loopLet = loopLet + 1" but set cannot have expression and also to reference a vector defined by let
  * we need to do "$&loopLet"
  let loopLet = $loopSet + 1 
  set loopSet = "$&loopLet"
  * to just change the device parameter use alter command
  * but to change the model paramater use altermod
  * also looks like spice is case insensitive hence M1 can also be written as m1
  altermod M1 lambda=$lmb
  echo #################################
  echo simulation for loopLet="$&loopLet" loopSet="$loopSet"
  * note this dc command is equivalent to the .dc inside the input deck, to execute the command inside the input deck use the run command
  DC Vds 0v 10v 100mv
  print V(1) I(Vds)
end

*let stop_r = 10k
*let delta_r = 1k
*let r_act = start_r
* loop
*while r_act le stop_r
*alter r1 r_act
*op
*print v(2)
*let r_act = r_act + delta_r
*end

echo Ending of control section
echo ++++++++++++++++++++++++++++++++++

.endc

.END

